//this will handle the timing restrictions aa required and stated in the user manual
//will be using the washer machine timer as a reference

//TS (Sync Pulse Time)
//  Vertical: Time- Clocks- Lines-
//  Horizontal: Time- Clocks-

//TDISP (Display Time)
//  Vertical: Time- Clocks- Lines-
//  Horizontal: Time- Clocks-

//TPW (Pulse Width)
//  Vertical: Time- Clocks- Lines-
//  Horizontal: Time- Clocks-

//TFP (Front Porch)
//  Vertical: Time- Clocks- Lines- 
//  Horizontal: Time- Clocks- 

//TBP (Back Porch)
//  Vertical: Time- Clocks- Lines-
//  Horizontal: Time- Clocks-

module vga_timer();

//Need to change names and values and erase Tw most likely

assign Ts = (counter >= );
   assign Tdisp =;
   assign Tpw =;
   assign Tfp = ;
   assign Tbp = ;

endmodule