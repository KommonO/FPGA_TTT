//Logic to handle the tic tac toe game for my final
//project in Rapid Prototyping with FPGAs
//Engineer: Kommon Ousley
//Date Started: 4/30/2016
//Inputs(May attempt to use the PS/2 Keyboard)
//
//Outputs
//player_1_win:1 bit wire
//player_2_win:1 bit wire
//
module ttt_logic(input mclk,  output wire player_1_win,player_2_win);

//wires
wire player1_turn, player2_turn;
wire enter;//also known as select depending on keyboard use or button use


//parameters
parameter 

	IDLE = ,	//IDLE state means that the screen is black
	START = ,	//Here we will also print the starting board 
	PLAYER1_MOVE = ,//takes in player 1's move, prints the new board, it is now player 2's turn
	PLAYER2_MOVE = ,//if it is player 2's turn in 



//logic block/state machine 1


//logic block/state machine 2




//clock process



//ASCII TEXT



endmodule
